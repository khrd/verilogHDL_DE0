module Lesson1(switch,led);

	inout switch;
	output led;
	
	assign led=switch;
	
endmodule